//  cw305_regs.vh
//  === Part of the side-channel measurement demo/proto.

`define REG_CLKSETTINGS     'h00
`define REG_USER_LED        'h01
`define REG_CRYPT_TYPE      'h02
`define REG_CRYPT_REV       'h03
`define REG_IDENTIFY        'h04
`define REG_TX_BYTE         'h05
`define REG_TX_IDX          'h06
`define REG_RX_BYTE         'h07
`define REG_RX_IDX          'h08
`define REG_RX_POS          'h09
`define REG_STATUS          'h0a
`define REG_BUILDTIME       'h0b

